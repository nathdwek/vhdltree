e1i1: entity e1
	e1i2 : entity e1
 e2I1:entity E2 --comment
E3i1:	entity lib.e3
