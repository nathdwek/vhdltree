chain: entity e5
