e1i1: entity long_component_name5678
	e1i2 : entity long_component_name5678
 e2I1:entity E2 --comment
E3_i1:	entity lib.e3
_badid: entity component
badid_: entity component
goodid1: entity .badcomponent
truncate_before_dot: entity e4.
bad_id_é"'(-è_ç)'": entity component
the: entity E_1
