on: entity e7
