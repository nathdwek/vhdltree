e3i2: entity lib.e3
