goes: entity e6
