long_ent17y_n4m3_with_numbers4567:  entity	lib.deep.E4
2numbers_should_not_start: entity component
