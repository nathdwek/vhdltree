--but stops
