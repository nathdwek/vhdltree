NO_PREFIX: entity e3
bad_prefix: entity lib.deep.e3
