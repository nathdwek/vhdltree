e4içàéè_éè_1:entity	lib.deep.E4
