check_recurse: entity lib.e3
NO_PREFIX: entity e3
bad_prefix: entity lib.deep.e3
